module controller(input wire 				clk,reset,
						input wire [31:12] 	Instr,
						input wire CO,N,Z,OVF,
						output wire 